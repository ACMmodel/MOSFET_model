** sch_path: /home/gmaranhao/Documents/MOSFET_model/Examples/GF180MCU/xschem/TB_not_acm.sch
**.subckt TB_not_acm
VA A VSS pulse(0 3.3 50n 200p 200p 50n 100n)
VDD VDD GND 3.3
VSS VSS GND 0
x1 A Y VDD VSS not_acm
**** begin user architecture code

.include /home/gmaranhao/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/gmaranhao/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.model NMOS_ACM nmos_ACM
.model PMOS_ACM pmos_ACM



.option gmin=1e-15

.control
pre_osdi ./NMOS_ACM_2V0.osdi
pre_osdi ./PMOS_ACM_2V0.osdi
save all


tran 1n 500n
remzerovec
write TB_not_acm.raw
set appendwrite

.endc


**** end user architecture code
**.ends

* expanding   symbol:  symbol/not_acm.sym # of pins=2
** sym_path: /home/gmaranhao/Documents/MOSFET_model/Examples/GF180MCU/xschem/symbol/not_acm.sym
** sch_path: /home/gmaranhao/Documents/MOSFET_model/Examples/GF180MCU/xschem/symbol/not_acm.sch
.subckt not_acm A Y VDDPIN VSSPIN
*.ipin A
*.opin Y
N1 Y A VSSPIN VSSPIN NMOS_ACM w=2u l=2u n=1.38 is=67.3n vt0=0.652 sigma=20m zeta=5m
N2 Y A VDDPIN VDDPIN PMOS_ACM w=2u l=2u n=1.438 is=17.94n vt0=0.7774 sigma=20m zeta=5m
.ends

.GLOBAL GND
.end
